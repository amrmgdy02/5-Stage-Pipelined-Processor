LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY ExecuteBlock IS
    PORT (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        ImmSignal : IN STD_LOGIC;
        InSignal : IN STD_LOGIC;
        InData : IN STD_LOGIC_VECTOR(15 DOWNTO 0); --data of in port
        Rs : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Source register 1
        Rt : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Source register 2
        WBEX_M : IN STD_LOGIC; -- Write-back enable from EX/MEM
        WBM_WB : IN STD_LOGIC; -- Write-back enable from MEM/WB
        RegDesE_M : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Destination register EX/MEM
        RegDesM_WB : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Destination register MEM/WB
        MemToReg_M_WB : IN STD_LOGIC; -- Memory-to-register signal from MEM/WB
        --Sel1FromForwarding : IN STD_LOGIC_VECTOR(1 DOWNTO 0); --ForwardA in forwarding unit
        --Sel2FromForwarding : IN STD_LOGIC_VECTOR(1 DOWNTO 0); --ForwardB in forwardingunit
        ReadData1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        ReadData2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        Immediate : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        AluSelector : IN STD_LOGIC_VECTOR(4 DOWNTO 0); --(basecode+opcode)
        AluResExecuteMemory : IN STD_LOGIC_VECTOR(15 DOWNTO 0); --Alu result which is stored in exexute memory register(alu to alu)
        WriteBackResult : IN STD_LOGIC_VECTOR(15 DOWNTO 0); --Same alu result but is stored in exexute memory writeback(memory to alu)
        -- ReadData1ExecuteMemory : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        -- ReadData1MemoryWriteBack : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       -- -MemOutMemoryWriteBack : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- it is the data output from memory
        --InPortExecuteMemory : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        --InPortMemoryWriteBack : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        ZeroFlag : OUT STD_LOGIC;
        NegativeFlag : OUT STD_LOGIC;
        CarryFlag : OUT STD_LOGIC;
        --OverflowFlag : OUT STD_LOGIC;
        AluOut : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- it is the data output from alu
        RsData : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- it is the data output from first upper mux 
        --ReadDataOut : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        --ReadDataOut2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        call_signal_in : IN STD_LOGIC;
        call_signal_out : OUT STD_LOGIC;
        save_flags : IN STD_LOGIC; -- Save current flags (INT)      --------------control signal to be added 
        rti_instruction_in : IN STD_LOGIC;
        restore_flags : IN STD_LOGIC; -- Restore saved flags (RTI)  --------------control signal to be added 
        restored_flags : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Flags to RESTORE FROM STACK
        --flags_out : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        update_flags : IN STD_LOGIC;
        --updated_flags : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        --ExecuteMemoryWriteBack : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        --conditional_branch : IN STD_LOGIC
        ------------------branching
        PCPlus1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Next sequential PC address
        ConditionalJumpZero : IN STD_LOGIC; -- Indicates a conditional jump (JZ)
        ConditionalJumpNegative : IN STD_LOGIC; -- Indicates a conditional jump (JN)
        ConditionalJumpCarry : IN STD_LOGIC; -- Indicates a conditional jump (JC)
        UnconditionalJump : IN STD_LOGIC; -- Indicates an unconditional jump (e.g., JMP, CALL, RET)
        FlushDecode : OUT STD_LOGIC;
        FlushExecute : OUT STD_LOGIC;
        ChangePC : OUT STD_LOGIC;
        NewPC : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        PCPlus1Out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0); --adddddddddddded
        rti_instruction_out : OUT STD_LOGIC;
		  store	: in std_logic
    );
    -- The updated_flags signal works alongside the update_flags control signal:
    -- If update_flags = '1', the execute block writes the new flags generated by the ALU (AluFlags).
    -- If update_flags = '0', the execute block passes the updated_flags value forward to preserve the existing flag state.
END ENTITY ExecuteBlock;

ARCHITECTURE Behavioral OF ExecuteBlock IS
    COMPONENT ALU IS
        GENERIC (n : INTEGER := 16);
        PORT (
            A, B : IN STD_LOGIC_VECTOR(n - 1 DOWNTO 0); -- Two operands
            Sel : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- Select lines
            FlagsIn : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Flags input (Zero, Negative,  Carry)
            FlagsOut : OUT STD_LOGIC_VECTOR(2 DOWNTO 0); -- Flags output (Zero, Negative,  Carry)
            Res : OUT STD_LOGIC_VECTOR(n - 1 DOWNTO 0) -- Result
            --BranchEnable : IN STD_LOGIC
        );
    END COMPONENT;

    COMPONENT FlagReg IS
        GENERIC (n : INTEGER := 3); -- Number of flags
        PORT (
            clk : IN STD_LOGIC; -- Clock signal
            rst : IN STD_LOGIC; -- Reset signal
            en : IN STD_LOGIC; -- Enable signal for writing flags
            flag : IN STD_LOGIC_VECTOR(n - 1 DOWNTO 0); -- Current flags to update (come from alu)
            flag_out : OUT STD_LOGIC_VECTOR(n - 1 DOWNTO 0); -- Output flags
            -- BranchEnable : IN STD_LOGIC; -- Clear Zero flag during branching
            save_flags : IN STD_LOGIC; -- Save current flags (INT)
            restore_flags : IN STD_LOGIC; -- Restore saved flags (RTI)
            restored_flags : IN STD_LOGIC_VECTOR(n - 1 DOWNTO 0); -- Flags to RESTORE FROM STACK
            saved_flags : OUT STD_LOGIC_VECTOR(n - 1 DOWNTO 0) -- Flags to save on interrupt
        );
    END COMPONENT;

    COMPONENT ForwardingUnit IS
        PORT (
            Rs : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Source register 1
            Rt : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Source register 2
            WBEX_M : IN STD_LOGIC; -- Write-back enable from EX/MEM
            WBM_WB : IN STD_LOGIC; -- Write-back enable from MEM/WB
            RegDesE_M : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Destination register EX/MEM
            RegDesM_WB : IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- Destination register MEM/WB
            MemToReg_M_WB : IN STD_LOGIC; -- Memory-to-register signal from MEM/WB
            ForwardA : OUT STD_LOGIC_VECTOR(1 DOWNTO 0); -- Forward control for ALU input A
            ForwardB : OUT STD_LOGIC_VECTOR(1 DOWNTO 0) -- Forward control for ALU input B
            ----UseMemResult : OUT STD_LOGIC -- Indicates if forwarding memory result
        );
    END COMPONENT;

    COMPONENT BranchingExecuteUnit IS
        PORT (
            reset : IN STD_LOGIC;
            ZeroFlag : IN STD_LOGIC; -- Flag for JZ (Jump if Zero)
            CarryFlag : IN STD_LOGIC; -- Flag for JC (Jump if Carry)
            NegativeFlag : IN STD_LOGIC; -- Flag for JN (Jump if Negative)
            PCPlus1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Next sequential PC address
            ConditionalJumpAddress : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- Address for conditional jumps
            ConditionalJumpZero : IN STD_LOGIC; -- Indicates a conditional jump (JZ)
            ConditionalJumpNegative : IN STD_LOGIC; -- Indicates a conditional jump (JN)
            ConditionalJumpCarry : IN STD_LOGIC; -- Indicates a conditional jump (JC)
            UnconditionalJump : IN STD_LOGIC; -- Indicates an unconditional jump (e.g., JMP, CALL, RET)
            FlushDecode : OUT STD_LOGIC; -- Control signal to flush the decode stage
            FlushExecute : OUT STD_LOGIC; -- Control signal to flush the execute stage
            ChangePC : OUT STD_LOGIC; -- Control signal to change the PC
            JumpAddress : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) -- Address to jump to
        );
    END COMPONENT;
    -- Internal signals
    SIGNAL Operand1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL Operand2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL Operand1_Final : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL Operand2_Final : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL Sel1FromForwarding : STD_LOGIC_VECTOR(1 DOWNTO 0);
    SIGNAL Sel2FromForwarding : STD_LOGIC_VECTOR(1 DOWNTO 0);
    SIGNAL AluResult : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL CurrentFlags : STD_LOGIC_VECTOR(2 DOWNTO 0); -- Current flags from Flag Register
    SIGNAL ALUFlagsOut : STD_LOGIC_VECTOR(2 DOWNTO 0); -- Flags output from ALU
    SIGNAL saved_flags : STD_LOGIC_VECTOR(2 DOWNTO 0); -- Flags saved in Flag Register
BEGIN
    -- Forwarding Unit instantiation
    ForwardingUnit_Instance : ForwardingUnit
    PORT MAP(
        Rs => Rs,
        Rt => Rt,
        WBEX_M => WBEX_M,
        WBM_WB => WBM_WB,
        RegDesE_M => RegDesE_M,
        RegDesM_WB => RegDesM_WB,
        MemToReg_M_WB => MemToReg_M_WB,
        ForwardA => Sel1FromForwarding,
        ForwardB => Sel2FromForwarding
    );
    -- Forwarding logic for Operand1
    PROCESS (Sel1FromForwarding, ReadData1, AluResExecuteMemory, WriteBackResult)
    BEGIN
        CASE Sel1FromForwarding IS
            WHEN "00" => Operand1 <= ReadData1;
            WHEN "01" => Operand1 <= AluResExecuteMemory;
            WHEN "10" => Operand1 <= WriteBackResult;
            WHEN OTHERS => Operand1 <= (OTHERS => '0');
        END CASE;
    END PROCESS;
    -- Forwarding logic for Operand2
    PROCESS (Sel2FromForwarding, ReadData2, AluResExecuteMemory, WriteBackResult)
    BEGIN
        -- forward a/b  --------> 00  ---->no forwarding
        --                        01  ---->Forward from EX/MEM
        --                        10  ---->Forward memory result from MEM/WB
        --                        11  ---->Forward ALU result from MEM/WB
        CASE Sel2FromForwarding IS
            WHEN "00" => Operand2 <= ReadData2;
            WHEN "01" => Operand2 <= AluResExecuteMemory;
            WHEN "10" => Operand2 <= WriteBackResult;
            WHEN OTHERS => Operand2 <= (OTHERS => '0');
        END CASE;

    END PROCESS;

    -- Logic to choose between Operand1 and InData based on InSignal
    PROCESS (InSignal, Operand1, InData)
    BEGIN
        IF InSignal = '1' THEN
            Operand1_Final <= InData; -- Use InData if InSignal is asserted
        ELSE
            Operand1_Final <= Operand1; -- Use Operand1 otherwise
        END IF;
    END PROCESS;

    -- Logic to choose between Operand2 and Immediate based on ImmSignal
    PROCESS (ImmSignal, Operand2, Immediate)
    BEGIN
        IF ImmSignal = '1' THEN
            Operand2_Final <= Immediate; -- Use Immediate if ImmSignal is asserted
        ELSE
            Operand2_Final <= Operand2; -- Use Operand2 otherwise
        END IF;
    END PROCESS;

    -- ALU instantiation
    ALU_Instance : ALU
    GENERIC MAP(n => 16)
    PORT MAP(
        A => Operand1_Final,
        B => Operand2_Final,
        Sel => AluSelector,
        FlagsIn => CurrentFlags, -- Flags from Flag Register
        FlagsOut => ALUFlagsOut, -- Flags output to Flag Register
        Res => AluResult
        --BranchEnable => call_signal_in
    );

    -- Flag Register instantiation
    FlagReg_Instance : FlagReg
    GENERIC MAP(n => 3)
    PORT MAP(
        clk => clk,
        rst => reset,
        en => update_flags, -- Enable signal to update flags
        flag => ALUFlagsOut, -- Flags from ALU
        flag_out => CurrentFlags, -- Current flags stored in register(i will take it and enter it as input in alu flags)
        save_flags => save_flags, -- Save flags signal during INTssss
        restore_flags => restore_flags, -- Restore flags signal during RTI
        restored_flags => restored_flags, -- Restore flags during RTI
        saved_flags => saved_flags -- Flags saved for interrupts (to be pushed in the stack)
    );

    BranchingUnit : BranchingExecuteUnit
    PORT MAP(
        reset => reset,
        ZeroFlag => ALUFlagsOut(0),
        CarryFlag => ALUFlagsOut(2),
        NegativeFlag => ALUFlagsOut(1),
        PCPlus1 => PCPlus1,
        ConditionalJumpAddress => AluResult,
        ConditionalJumpZero => ConditionalJumpZero,
        ConditionalJumpNegative => ConditionalJumpNegative,
        ConditionalJumpCarry => ConditionalJumpCarry,
        UnconditionalJump => UnconditionalJump,
        FlushDecode => FlushDecode,
        FlushExecute => FlushExecute,
        ChangePC => ChangePC,
        JumpAddress => NewPC
    );

    RsData <= Operand1 when store ='0' else Operand2;
    AluOut <= AluResult;
    ZeroFlag <= CurrentFlags(0);
    NegativeFlag <= CurrentFlags(1);
    CarryFlag <= CurrentFlags(2);
    PCPlus1Out <= saved_flags & PCPlus1(12 DOWNTO 0); -------added now flags stored in last 3 bits 
    rti_instruction_out <= rti_instruction_in;
    call_signal_out <= call_signal_in;

END ARCHITECTURE Behavioral;